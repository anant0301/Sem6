`include"and64_16.v"
module and64_32(
	input [63:0] in1,
	input [31:0] in2,
	output [63:0] out0,
	output [63:0] out1,
	output [63:0] out2,
	output [63:0] out3,
	output [63:0] out4,
	output [63:0] out5,
	output [63:0] out6,
	output [63:0] out7,
	output [63:0] out8,
	output [63:0] out9,
	output [63:0] out10,
	output [63:0] out11,
	output [63:0] out12,
	output [63:0] out13,
	output [63:0] out14,
	output [63:0] out15,
	output [63:0] out16,
	output [63:0] out17,
	output [63:0] out18,
	output [63:0] out19,
	output [63:0] out20,
	output [63:0] out21,
	output [63:0] out22,
	output [63:0] out23,
	output [63:0] out24,
	output [63:0] out25,
	output [63:0] out26,
	output [63:0] out27,
	output [63:0] out28,
	output [63:0] out29,
	output [63:0] out30,
	output [63:0] out31
);
	and64_16 a0(
		in1[63:0], 
		in2[15:0], 
		out0[63:0],
		out1[63:0],
		out2[63:0],
		out3[63:0],
		out4[63:0],
		out5[63:0],
		out6[63:0],
		out7[63:0],
		out8[63:0],
		out9[63:0],
		out10[63:0],
		out11[63:0],
		out12[63:0],
		out13[63:0],
		out14[63:0],
		out15[63:0]
		);
	and64_16 a1(
		in1[63:0], 
		in2[31:16], 
		out16[63:0],
		out17[63:0],
		out18[63:0],
		out19[63:0],
		out20[63:0],
		out21[63:0],
		out22[63:0],
		out23[63:0],
		out24[63:0],
		out25[63:0],
		out26[63:0],
		out27[63:0],
		out28[63:0],
		out29[63:0],
		out30[63:0],
		out31[63:0]
		);
endmodule

